CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
40 0 6 110 10
176 80 1364 747
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
76546066 0
0
6 Title:
5 Name:
0
0
0
10
2 +V
167 294 256 0 1 3
0 14
0
0 0 54256 0
2 5V
-7 -22 7 -14
2 V2
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
762 0 0
2
5.89883e-315 0
0
7 Pulser~
4 206 408 0 10 12
0 17 18 12 19 0 0 5 5 1
7
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
39 0 0
2
5.89883e-315 0
0
9 CC 7-Seg~
183 947 178 0 18 19
10 8 7 6 5 4 3 2 20 21
0 0 0 1 1 1 1 2 2
0
0 0 21088 0
6 BLUECC
13 -41 55 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
9450 0 0
2
5.89883e-315 0
0
9 2-In AND~
219 685 230 0 3 22
0 15 13 16
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
3236 0 0
2
5.89883e-315 0
0
9 2-In AND~
219 523 222 0 3 22
0 10 9 15
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
3321 0 0
2
5.89883e-315 0
0
6 74112~
219 757 335 0 7 32
0 14 16 12 16 14 22 11
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U3B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 2 0
1 U
8879 0 0
2
5.89883e-315 0
0
6 74112~
219 610 333 0 7 32
0 14 15 12 15 14 13 13
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U3A
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 0 2 1 2 0
1 U
5433 0 0
2
5.89883e-315 0
0
6 74112~
219 441 336 0 7 32
0 14 10 12 10 14 23 9
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U2B
22 -61 43 -53
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 10 11 13 12 14 7 9 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 1 0
1 U
3679 0 0
2
5.89883e-315 0
0
6 74112~
219 294 336 0 7 32
0 14 14 12 14 14 24 10
0
0 0 4720 0
5 74112
4 -60 39 -52
3 U2A
21 -62 42 -54
0
15 DVCC=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 4 3 1 2 15 6 5 4 3
1 2 15 6 5 10 11 13 12 14
7 9 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 1 0
1 U
9342 0 0
2
5.89883e-315 0
0
6 74LS48
188 910 353 0 14 29
0 11 13 9 10 25 26 2 3 4
5 6 7 8 27
0
0 0 4848 90
6 74LS48
-21 -60 21 -52
2 U1
57 -3 71 5
0
15 DVCC=16;DGND=8;
119 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %14i]
+ [%16bo %1o %2o %3o %4o %5o %6o %14o %7o %8o %9o %10o %11o %12o %13o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 3 5 14 15 9
10 11 12 13 4 6 2 1 7 3
5 14 15 9 10 11 12 13 4 0
65 0 0 512 1 0 0 0
1 U
3623 0 0
2
5.89883e-315 0
0
36
7 7 2 0 0 12416 0 10 3 0 0 4
872 323
872 305
962 305
962 214
8 6 3 0 0 12416 0 10 3 0 0 4
881 323
881 296
956 296
956 214
9 5 4 0 0 12416 0 10 3 0 0 4
890 323
890 287
950 287
950 214
10 4 5 0 0 12416 0 10 3 0 0 4
899 323
899 279
944 279
944 214
11 3 6 0 0 12416 0 10 3 0 0 4
908 323
908 272
938 272
938 214
12 2 7 0 0 4224 0 10 3 0 0 4
917 323
917 265
932 265
932 214
13 1 8 0 0 4224 0 10 3 0 0 2
926 323
926 214
0 3 9 0 0 8320 0 0 10 26 0 4
492 300
492 425
890 425
890 387
0 4 10 0 0 8320 0 0 10 36 0 4
333 300
333 438
899 438
899 387
7 1 11 0 0 8320 0 6 10 0 0 5
781 299
824 299
824 401
872 401
872 387
3 0 12 0 0 4096 0 2 0 0 33 2
230 399
260 399
6 0 13 0 0 4096 0 7 0 0 13 2
640 315
652 315
0 2 13 0 0 16512 0 0 10 28 0 6
652 297
652 315
683 315
683 414
881 414
881 387
0 1 14 0 0 8192 0 0 1 23 0 4
243 300
243 266
294 266
294 265
1 0 14 0 0 0 0 1 0 0 19 2
294 265
294 265
0 0 14 0 0 4096 0 0 0 19 22 2
355 265
355 356
1 1 14 0 0 8192 0 7 6 0 0 4
610 270
610 265
757 265
757 272
1 1 14 0 0 8320 0 8 7 0 0 4
441 273
441 265
610 265
610 270
1 1 14 0 0 0 0 9 8 0 0 4
294 273
294 265
441 265
441 273
5 5 14 0 0 0 0 7 6 0 0 4
610 345
610 356
757 356
757 347
5 5 14 0 0 0 0 8 7 0 0 4
441 348
441 356
610 356
610 345
5 5 14 0 0 0 0 9 8 0 0 4
294 348
294 356
441 356
441 348
4 2 14 0 0 0 0 9 9 0 0 4
270 318
243 318
243 300
270 300
2 0 15 0 0 4096 0 7 0 0 25 2
586 297
548 297
0 4 15 0 0 4224 0 0 7 27 0 3
548 221
548 315
586 315
2 7 9 0 0 0 0 5 8 0 0 4
499 231
492 231
492 300
465 300
3 1 15 0 0 12416 0 5 4 0 0 4
544 222
548 222
548 221
661 221
2 7 13 0 0 0 0 4 7 0 0 4
661 239
652 239
652 297
634 297
2 0 16 0 0 4096 0 6 0 0 30 2
733 299
712 299
3 4 16 0 0 8320 0 4 6 0 0 4
706 230
712 230
712 317
733 317
3 0 12 0 0 8192 0 7 0 0 33 3
580 306
576 306
576 399
3 0 12 0 0 0 0 8 0 0 33 3
411 309
405 309
405 399
3 3 12 0 0 12432 0 9 6 0 0 6
264 309
260 309
260 399
725 399
725 308
727 308
1 0 10 0 0 0 0 5 0 0 35 3
499 213
383 213
383 300
4 0 10 0 0 0 0 8 0 0 36 3
417 318
383 318
383 300
7 2 10 0 0 0 0 9 8 0 0 2
318 300
417 300
1
-16 0 0 0 400 0 0 0 0 3 2 1 34
14 Century Gothic
0 0 0 35
404 79 742 104
413 86 732 105
35 BINARY 4-BIT SYNCHRONOUS UP COUNTER
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
